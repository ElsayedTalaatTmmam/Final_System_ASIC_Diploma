
`timescale 1ns/1ps

module SYS_TOP_TB ();

/////////////////////////////////////////////////////////
///////////////////// Parameters ////////////////////////
/////////////////////////////////////////////////////////

parameter DATA_WIDTH_TB  = 8  ;
parameter ADDR_WIDTH_TB  = 4  ;   
parameter REF_CLK_PER = 10 ;         // 100 MHz
parameter UART_CLK_PER = 271.267 ;   // 3.6864 MHz (115.2 * 32)

parameter WR_CMD  = 8'hAA ;          // write coomand
parameter RD_CMD  = 8'hBB ;          // read command  
parameter ALU_WOP_CMD  = 8'hCC ;     // write operation ( from TB ) 
parameter ALU_WNOP_CMD = 8'hDD ;     // write 

/////////////////////////////////////////////////////////
//////////////////// DUT Signals ////////////////////////
/////////////////////////////////////////////////////////

reg                                RST_N;
reg                                UART_CLK;
reg                                REF_CLK;
reg                                UART_RX_IN;
wire                               UART_TX_O;
wire                               parity_error;
wire                               framing_error;

////////////////////////////////////////////////////////
////////////////// initial block /////////////////////// 
////////////////////////////////////////////////////////

initial
 begin

 // Initialization
 initialize() ;
 // Reset
 reset() ; 

 ////////////////   Configuration 1     //////////////////
 ////////////////   PRESCALE : 32       //////////////////
 ////////////////   Parity   : Enabled  //////////////////
 ////////////////   TYPE     : EVEN     //////////////////
   SEND_WR_CMD(8'h02,8'h81) ;
 //SEND_WR_CMD(8'h02,8'h81) ;

 /////////////////////  WRITE CMD  ///////////////////////
  //Send Write Command (Address:8'h06 & Data: 8'hA5)
  SEND_WR_CMD(8'h06,8'hA5) ;
 
  //Check Write Operation
  CHECK_WR(8'h06,8'hA5) ;

 /////////////////////  READ CMD   ///////////////////////
  // Send Read Command (Address:8'h02)
  SEND_RD_CMD(8'h02) ;
 
  // Check Read Operation
  CHECK_RD(8'h02) ;

 ////////////////////  ALU_WOP CMD   ////////////////////
  // Send ALU WOP Command (OP_A = 100 & OP_B = 50 & FUNC = Subtraction)
$display ("//*********************** ALU Operation A/B from INPUT ********************************//");
  SEND_ALU_WOP_CMD(8'd100,8'd50,8'd1) ;

  // Check ALU Command
  CHECK_ALU(8'd1) ;
 //////////////////// ALU_WNOP CMD //////////////////////
  // Send ALU WNOP Command (FUNC = Addition)
$display ("//*********************** ALU Operation A/B from RAM **********************************//");
  SEND_ALU_WNOP_CMD(8'd1) ;

  // Check ALU Command
  CHECK_ALU(8'd1) ;
                        $display(" << ---------------------------------------------------------------------------------------- >>");

 ///////////////////////////////////////////////////////// 
 ////////////////   Configuration 2     //////////////////
 ////////////////   PRESCALE : 32       //////////////////
 ////////////////   Parity   : Enabled  //////////////////
 ////////////////   TYPE     : ODD      ////////////////// 
 /////////////////////////////////////////////////////////

 SEND_WR_CMD(8'h02,8'h83) ;

 /////////////////////  WRITE CMD  ///////////////////////
  //Send Write Command (Address:8'h06 & Data: 8'hA5)
  SEND_WR_CMD(8'h0A,8'h19) ;
 
  //Check Write Operation
  CHECK_WR(8'h0A,8'h19) ;

 /////////////////////  READ CMD   ///////////////////////
  // Send Read Command (Address:8'h02)
  SEND_RD_CMD(8'h02) ;
 
  // Check Read Operation
  CHECK_RD(8'h02) ;

 ////////////////////  ALU_WOP CMD   ////////////////////
  // Send ALU WOP Command (OP_A = 100 & OP_B = 50 & FUNC = Subtraction)
$display ("//*********************** ALU Operation A/B from INPUT ********************************//");
  SEND_ALU_WOP_CMD(8'd120,8'd80,8'd1) ;
  // Check ALU Command
  CHECK_ALU(8'd1) ;

 //////////////////// ALU_WNOP CMD //////////////////////
  // Send ALU WNOP Command (FUNC = Addition)
$display ("//*********************** ALU Operation A/B from RAM **********************************//");
  SEND_ALU_WNOP_CMD(8'd0) ;
 
  // Check ALU Command
  CHECK_ALU(8'd0) ;  
                        $display(" << ---------------------------------------------------------------------------------------- >>");

 ///////////////////////////////////////////////////////// 
 ////////////////   Configuration 3     //////////////////
 ////////////////   PRESCALE : 32       //////////////////
 ////////////////   Parity   : DISABLED //////////////////
 /////////////////////////////////////////////////////////

 SEND_WR_CMD(8'h02,8'h80) ;

 /////////////////////  WRITE CMD  ///////////////////////
  //Send Write Command (Address:8'h06 & Data: 8'hA5)
  SEND_WR_CMD(8'h08,8'h75) ;
 
  //Check Write Operation
  CHECK_WR(8'h08,8'h75) ;

 /////////////////////  READ CMD   ///////////////////////
  // Send Read Command (Address:8'h02)
  SEND_RD_CMD(8'h06) ;
 
  // Check Read Operation
  CHECK_RD(8'h06) ;

 ////////////////////  ALU_WOP CMD   ////////////////////
  // Send ALU WOP Command (OP_A = 100 & OP_B = 50 & FUNC = Subtraction)
$display ("//*********************** ALU Operation A/B from INPUT ********************************//");
  SEND_ALU_WOP_CMD(8'd100,8'd50,8'd1) ;
 
  // Check ALU Command
  CHECK_ALU(8'd1) ;

 //////////////////// ALU_WNOP CMD //////////////////////
  // Send ALU WNOP Command (FUNC = Addition)
$display ("//*********************** ALU Operation A/B from RAM **********************************//");
  SEND_ALU_WNOP_CMD(8'd0) ;
 
  // Check ALU Command
  CHECK_ALU(8'd0) ;  
                        $display(" << ---------------------------------------------------------------------------------------- >>");

#400
$stop ;
end

////////////////////////////////////////////////////////
/////////////////////// TASKS //////////////////////////
////////////////////////////////////////////////////////

/////////////// Signals Initialization //////////////////

task initialize ;
  begin
	UART_CLK          = 1'b0   ;
	REF_CLK           = 1'b0   ;
	RST_N             = 1'b1   ;    // rst is deactivated
	UART_RX_IN        = 1'b1   ;
  end
endtask

///////////////////////// RESET /////////////////////////
task reset ;
  begin
	#(REF_CLK_PER)
	RST_N  = 'b0;           // rst is activated
	#(REF_CLK_PER)
	RST_N  = 'b1;
	#(REF_CLK_PER) ;
  end
endtask

/////////////////////// Load Frame /////////////////////////   /****  strt -- data -- parity -- stop  ****/

task LD_FRAME ;
   input  [DATA_WIDTH_TB-1:0]  FRAME_DATA ;
   integer   i  ; 
 begin
      @ (posedge DUT.UART_TX_U0.CLK)  
	UART_RX_IN <= 1'b0 ;                    // start_bit
	for(i=0; i<8; i=i+1)
		begin
		@(posedge DUT.UART_TX_U0.CLK) 		
		UART_RX_IN <= FRAME_DATA[i] ;       // frame data bits
		end 

	if(DUT.U0_RegFile.REG2[0])                               /// if Enable 
		begin                                            /* calculate PARITY bit */
			@ (posedge DUT.UART_TX_U0.CLK) 
			case(DUT.U0_RegFile.REG2[1])
			1'b0 : UART_RX_IN <= ^FRAME_DATA  ;     // Even Parity
			1'b1 : UART_RX_IN <= ~^FRAME_DATA ;     // Odd Parity
			endcase	
		end
	@ (posedge DUT.UART_TX_U0.CLK) 
	UART_RX_IN <= 1'b1 ;              // stop_bit	
 end
endtask 

/////////////////////// WRITE CMD /////////////////////////
task SEND_WR_CMD ;
  input  [DATA_WIDTH_TB-1:0]  ADDR ;
  input  [DATA_WIDTH_TB-1:0]  DATA ;
 begin
	LD_FRAME(WR_CMD) ;   // Load Write Command
	LD_FRAME(ADDR)   ;   // Load Write Address
	LD_FRAME(DATA)	 ;   // Load Write Data
 end
endtask 

/////////////////////// Read CMD /////////////////////////
task SEND_RD_CMD ;
    input  [DATA_WIDTH_TB-1:0]  ADDR ;
 begin
	LD_FRAME(RD_CMD) ;  // Load Read Command
	LD_FRAME(ADDR)   ;  // Load Read Address
 end
endtask 

///////////////////// ALU_WOP CMD ///////////////////////
task SEND_ALU_WOP_CMD ;
   input  [DATA_WIDTH_TB-1:0]  OP_A ;
   input  [DATA_WIDTH_TB-1:0]  OP_B ;
   input  [DATA_WIDTH_TB-1:0]  FUNC ;
 begin
	LD_FRAME(ALU_WOP_CMD) ;	   // Load ALU_WOP Command
	LD_FRAME(OP_A)        ;    // Load Operand A 
	LD_FRAME(OP_B)	      ;    // Load Operand B 
	LD_FRAME(FUNC)        ;    // Load ALU Function
 end
endtask 

///////////////////// ALU_WOP CMD ///////////////////////
task SEND_ALU_WNOP_CMD ;
   input  [DATA_WIDTH_TB-1:0]  FUNC ; 
 begin
	LD_FRAME(ALU_WNOP_CMD)	 ;    // Load ALU_WOP Command
	LD_FRAME(FUNC)           ;    // Load ALU Function
 end
endtask 

//////////////// Check Write Operation /////////////////
task CHECK_WR ;
   input  [DATA_WIDTH_TB-1:0]  ADDR ;
   input  [DATA_WIDTH_TB-1:0]  DATA ; 
 begin
	wait(DUT.U0_RegFile.WrEn)              // after SYS_CTRL WrEn =1
	repeat(2) @(posedge REF_CLK); 
	if(DUT.U0_RegFile.memory[ADDR[ADDR_WIDTH_TB-1:0]] == DATA)
		begin
			$display("Write Operation is succeeded / PARITY_EN=%d PARITY_TYPE=%d  PRESCALE=%d  ",DUT.U0_RegFile.REG2[0],DUT.U0_RegFile.REG2[1],DUT.U0_RegFile.REG2[7:2]);
		end
	else
		begin
			$display("Write Operation is failed / PARITY_EN=%d PARITY_TYPE=%d  PRESCALE=%d  ",DUT.U0_RegFile.REG2[0],DUT.U0_RegFile.REG2[1],DUT.U0_RegFile.REG2[7:2]);
		end	
 end
endtask 

//////////////// Check Read Operation /////////////////
task CHECK_RD ;
  input  [DATA_WIDTH_TB-1:0]  	ADDR     ; 
     reg    [10:0]  gener_out ,expec_out;     //longest frame = 11 bits (1-start,1-stop,8-data,1-parity)
     reg            parity_bit;
   integer   i  ;
 begin
	//generated frame
	@(posedge DUT.UART_TX_U0.busy)                                  // after load data at UART_TX
	for(i=0; i<11; i=i+1)
		begin
		@(negedge DUT.UART_TX_U0.CLK) gener_out[i] = UART_TX_O ;
		end	
	//calculate expected parity bit 	
    if(DUT.U0_RegFile.REG2[0])
		if(DUT.U0_RegFile.REG2[1])
			parity_bit = ~^DUT.U0_RegFile.memory[ADDR[ADDR_WIDTH_TB-1:0]] ;
		else
			parity_bit = ^DUT.U0_RegFile.memory[ADDR[ADDR_WIDTH_TB-1:0]] ;
         	else
			parity_bit = 1'b1 ;		
	//expected frame
    if(DUT.U0_RegFile.REG2[0])
		expec_out = {1'b1,parity_bit,DUT.U0_RegFile.memory[ADDR[ADDR_WIDTH_TB-1:0]],1'b0} ;
	else
		expec_out = {1'b1,1'b1,DUT.U0_RegFile.memory[ADDR[ADDR_WIDTH_TB-1:0]],1'b0} ;
			
	if(gener_out == expec_out) 
		begin
			$display(" Read Operation is succeeded / PARITY_EN=%d PARITY_TYPE=%d  PRESCALE=%d  ",DUT.U0_RegFile.REG2[0],DUT.U0_RegFile.REG2[1],DUT.U0_RegFile.REG2[7:2]);
		end
	else
		begin
			$display(" Read Operation is failed / PARITY_EN=%d PARITY_TYPE=%d  PRESCALE=%d  ",DUT.U0_RegFile.REG2[0],DUT.U0_RegFile.REG2[1],DUT.U0_RegFile.REG2[7:2]);
		end
 end
endtask

//////////////// Check ALU Operation /////////////////
task CHECK_ALU ;
  input  [DATA_WIDTH_TB-1:0]  	FUNCTION ;
 //longest frame = 11 bits (1-start,1-stop,8-data,1-parity) 
   reg    [10:0]  gener_byte0  , gener_byte1 ;     
   reg    [10:0]  expec_byte0  , expec_byte1  ;                        
   reg            parity_bit0 , parity_bit1 ; 
   reg    [2*DATA_WIDTH_TB-1:0] ALU_OUT_RESULT ; 
     integer   i  ;
 begin
	//generated byte0 frame
	@(posedge DUT.UART_TX_U0.busy)                  // first byte 
	for(i=0; i<11; i=i+1)
		begin
		@(negedge DUT.UART_TX_U0.CLK) gener_byte0[i] = UART_TX_O ;
		end		

	//generated byte1 frame
	@(posedge DUT.UART_TX_U0.busy)                   // second byte 
	for(i=0; i<11; i=i+1)
		begin
		@(negedge DUT.UART_TX_U0.CLK) gener_byte1[i] = UART_TX_O ;

		end		
	//calculate ALU Output  	
	case (FUNCTION) 
     4'b0000: begin   ALU_OUT_RESULT = DUT.U0_RegFile.memory[0] + DUT.U0_RegFile.memory[1];              end
     4'b0001: begin   ALU_OUT_RESULT = DUT.U0_RegFile.memory[0] - DUT.U0_RegFile.memory[1];              end
     4'b0010: begin   ALU_OUT_RESULT = DUT.U0_RegFile.memory[0] * DUT.U0_RegFile.memory[1];              end
     4'b0011: begin   ALU_OUT_RESULT = DUT.U0_RegFile.memory[0] / DUT.U0_RegFile.memory[1];              end
     4'b0100: begin   ALU_OUT_RESULT = DUT.U0_RegFile.memory[0] & DUT.U0_RegFile.memory[1];              end
     4'b0101: begin   ALU_OUT_RESULT = DUT.U0_RegFile.memory[0] | DUT.U0_RegFile.memory[1];              end
     4'b0110: begin   ALU_OUT_RESULT = ~ (DUT.U0_RegFile.memory[0] & DUT.U0_RegFile.memory[1]);          end
     4'b0111: begin   ALU_OUT_RESULT = ~ (DUT.U0_RegFile.memory[0] | DUT.U0_RegFile.memory[1]);          end     
     4'b1000: begin   ALU_OUT_RESULT =  (DUT.U0_RegFile.memory[0] ^ DUT.U0_RegFile.memory[1]);           end
     4'b1001: begin   ALU_OUT_RESULT = ~ (DUT.U0_RegFile.memory[0] ^ DUT.U0_RegFile.memory[1]);          end           
     4'b1010: begin
              if (DUT.U0_RegFile.memory[0] == DUT.U0_RegFile.memory[1])     ALU_OUT_RESULT = 'b1;
              else                                                          ALU_OUT_RESULT = 'b0;        end
     4'b1011: begin
               if (DUT.U0_RegFile.memory[0] > DUT.U0_RegFile.memory[1])     ALU_OUT_RESULT = 'b10;
               else                                                         ALU_OUT_RESULT = 'b0;        end 
     4'b1100: begin
               if (DUT.U0_RegFile.memory[0] < DUT.U0_RegFile.memory[1])     ALU_OUT_RESULT = 'b11;
               else                                                         ALU_OUT_RESULT = 'b0;        end     
     4'b1101: begin               ALU_OUT_RESULT = DUT.U0_RegFile.memory[0]>>1;                          end
     4'b1110: begin               ALU_OUT_RESULT = DUT.U0_RegFile.memory[0]<<1;                          end
     4'b1111: begin               ALU_OUT_RESULT = 'b0;                                                  end
    endcase

	//calculate expected parity bit for ALU byte0 data  	
    if(DUT.U0_RegFile.REG2[0])
		if(DUT.U0_RegFile.REG2[1])    parity_bit0 = ~^ALU_OUT_RESULT[DATA_WIDTH_TB-1:0] ;
		else        		      parity_bit0 = ^ALU_OUT_RESULT[DATA_WIDTH_TB-1:0] ;
	else        parity_bit0 = 1'b1 ;	

	//calculate expected parity bit for ALU byte1 data  	
    if(DUT.U0_RegFile.REG2[0])
		if(DUT.U0_RegFile.REG2[1])    parity_bit1 = ~^ALU_OUT_RESULT[2*DATA_WIDTH_TB-1:DATA_WIDTH_TB] ;
		else   			      parity_bit1 = ^ALU_OUT_RESULT[2*DATA_WIDTH_TB-1:DATA_WIDTH_TB] ;
	else        parity_bit1 = 1'b1 ;	

	//expected byte0 frame 
    if(DUT.U0_RegFile.REG2[0])		expec_byte0 = {1'b1,parity_bit0,ALU_OUT_RESULT[DATA_WIDTH_TB-1:0],1'b0} ;
	else            		expec_byte0 = {1'b1,1'b1,ALU_OUT_RESULT[DATA_WIDTH_TB-1:0],1'b0} ;

	//expected byte1 frame 
    if(DUT.U0_RegFile.REG2[0])		expec_byte1 = {1'b1,parity_bit1,ALU_OUT_RESULT[2*DATA_WIDTH_TB-1:DATA_WIDTH_TB],1'b0} ;
	else            		expec_byte1 = {1'b1,1'b1,ALU_OUT_RESULT[2*DATA_WIDTH_TB-1:DATA_WIDTH_TB],1'b0} ;

	if(gener_byte0 == expec_byte0 && gener_byte1 == expec_byte1) 
		begin
			$display("  ALU Operation is succeeded / PARITY_EN=%d PARITY_TYPE=%d  PRESCALE=%d  ",DUT.U0_RegFile.REG2[0],DUT.U0_RegFile.REG2[1],DUT.U0_RegFile.REG2[7:2]);
		end
	else
		begin
			$display("  ALU Operation is failed / PARITY_EN=%d PARITY_TYPE=%d  PRESCALE=%d  ",DUT.U0_RegFile.REG2[0],DUT.U0_RegFile.REG2[1],DUT.U0_RegFile.REG2[7:2]);
                end
	end
endtask

//////////////////////////////////////////////////////// 
///////////////////// Clock Generator //////////////////
////////////////////////////////////////////////////////
 
// REF Clock Generator
always #(REF_CLK_PER/2) REF_CLK = ~REF_CLK ;

// UART RX Clock Generator
always #(UART_CLK_PER/2) UART_CLK = ~UART_CLK ;

//////////////////////////////////////////////////////// 
///////////////// Design Instaniation //////////////////
////////////////////////////////////////////////////////

SYS_TOP # (.DATA_WIDTH(DATA_WIDTH_TB) ,  .RF_ADDR(ADDR_WIDTH_TB)) DUT (
.UART_CLK(UART_CLK),
.REF_CLK(REF_CLK),
.RST_N(RST_N),
.UART_RX_IN(UART_RX_IN),
.UART_TX_O(UART_TX_O),
.parity_error(parity_error),
.framing_error(framing_error)
);

endmodule 